library verilog;
use verilog.vl_types.all;
entity UpDownBinaryCounter_vlg_vec_tst is
end UpDownBinaryCounter_vlg_vec_tst;
