library verilog;
use verilog.vl_types.all;
entity nandgate_vlg_vec_tst is
end nandgate_vlg_vec_tst;
