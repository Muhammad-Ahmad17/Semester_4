library verilog;
use verilog.vl_types.all;
entity FourBitCounter_vlg_vec_tst is
end FourBitCounter_vlg_vec_tst;
